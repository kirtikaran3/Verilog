`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   13:17:57 02/08/2017
// Design Name:   ortest
// Module Name:   C:/Users/Kirti/Documents/verilog/PTUVLSI/andTest/ortb.v
// Project Name:  andTest
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ortest
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module ortb;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	ortest uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

