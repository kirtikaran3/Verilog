$date
   Sat Jan 28 12:05:46 2017
$end
$version
  P.28xd
$end
$timescale
  1ps
$end
$scope module tb $end
$var wire 1 & out $end
$var reg 1 " a $end
$var reg 1 # b $end
$scope module uut $end
$var wire 1 $ a $end
$var wire 1 % b $end
$var wire 1 & out $end
$upscope $end
$upscope $end
$enddefinitions $end
#100000
$dumpvars
0"
0#
0$
0%
0&
$end
#110000
1#
1%
#115000
1"
0#
1$
0%
#120000
1#
$dumpoff
x&
x$
x%
x&
x"
x#
$end
