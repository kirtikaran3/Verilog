`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:29:22 11/15/2016 
// Design Name: 
// Module Name:    andgatetest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module andgatetest(in0,in1,out    );

	input in0,in1; 
	output out; 
	
	assign out = in0 & in1;


endmodule





