`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:27:46 01/21/2017 
// Design Name: 
// Module Name:    ass 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ass(
   in,out,clk );


input in,clk; 
output out; 
reg out; 

always @(posedge clk) 
begin 

		 out = in;

end 


endmodule









