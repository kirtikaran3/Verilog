`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:16:28 04/14/2016 
// Design Name: 
// Module Name:    assdeass 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module assdeass(in,out,clk    );

input in,clk; 
output out; 
reg out; 

always @(posedge clk) 

	begin 

	assign	 out=in;

	end


endmodule





















