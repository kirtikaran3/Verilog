`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:26:30 01/28/2017 
// Design Name: 
// Module Name:    andUDP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module andUDP(
 a,b,o   );

input a,b; 
output o; 

new

new(o,a,b);
 

endmodule

primitive new(o,a,b); 

output o; 
input a,b; 

table  

	0	0:	0; 
	1	0:	0; 
	0	1:	0; 
	1	1:	1;


endtable 




endprimitive


